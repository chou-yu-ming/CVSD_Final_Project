package dat_0;
integer pat_num = 0;
reg [767:0] input_data  = 768'h259f4329e6f4590b9a164106cf6a659eb4862b21fb97d43588561712e8e5216a0fa4d2a95dafe3275eaf3ba907dbb1da819aba3927450d7399a270ce660d2fae2f0fe2678dedf6671e055f1a557233b324f44fb8be4afe607e5541eb11b0bea2;
reg [511:0] golden_data = 512'h47f6a5d15e1a09495f9216eba5253538db62c06ad333adbcc86932c069f00d26465032bc1d1cace745d1b3bad5ca1115805ab1512361151d1c84c68aa2f54468;
endpackage

package dat_1;
integer pat_num = 1;
reg [767:0] input_data  = 768'h17e0aa3c03983ca8ea7e9d498c778ea6eb2083e6ce164dba0ff18e0242af9fc32e2c9fbf00b87ab7cde15119d1c5b09aa9743b5c6fb96ec59dbf2f30209b133c116943db82ba4a31f240994b14a091fb55cc6edd19658a06d5f4c5805730c232;
reg [511:0] golden_data = 512'h7a3afed80c2ab24733d7a3cf8b33efcd547e88fabc71b39da58b42a26e6c606c6cbfdc595891983cc17335e1ecfbd786b92805efbd5be956a142f23285f29f8c;
endpackage

package dat_2;
integer pat_num = 2;
reg [767:0] input_data  = 768'h1759edc372ae22448b0163c1cd9d2b7d247a8333f7b0b7d2cda8056c3d15eef75b90ea17eaf962ef96588677a54b09c016ad982c842efa107c078796f88449a86a210d43f514ec3c7a8e677567ad835b5c2e4bc5dd3480e135708e41b42c0ac6;
reg [511:0] golden_data = 512'h668e7ea762ae11fb5159d50df7f92ee488c0f5ac4266701687de38e61cc5c8062bc1a2c8137938914f9b6e42763026845c6ee2c134819c7ba755a513d05c6ec8;
endpackage